-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Sat May 27 10:11:26 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY stateMachineDec IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        aceptar : IN STD_LOGIC := '0';
        Q1 : OUT STD_LOGIC;
        Q0 : OUT STD_LOGIC;
        letra0 : OUT STD_LOGIC;
        letra1 : OUT STD_LOGIC;
        letra2 : OUT STD_LOGIC;
        letra3 : OUT STD_LOGIC
    );
END stateMachineDec;

ARCHITECTURE BEHAVIOR OF stateMachineDec IS
    TYPE type_fstate IS (ptosGanar,avisoRonda,inputRonda,ptosJugadores,registroPtos,inputPtos);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,aceptar)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= ptosGanar;
            Q1 <= '0';
            Q0 <= '0';
            letra0 <= '0';
            letra1 <= '0';
            letra2 <= '0';
            letra3 <= '0';
        ELSE
            Q1 <= '0';
            Q0 <= '0';
            letra0 <= '0';
            letra1 <= '0';
            letra2 <= '0';
            letra3 <= '0';
            CASE fstate IS
                WHEN ptosGanar =>
                    IF ((aceptar = '1')) THEN
                        reg_fstate <= avisoRonda;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ptosGanar;
                    END IF;

                    letra3 <= '1';

                    letra2 <= '1';

                    letra1 <= '1';

                    letra0 <= '0';

                    Q0 <= '1';

                    Q1 <= '0';
                WHEN avisoRonda =>
                    IF ((aceptar = '1')) THEN
                        reg_fstate <= inputRonda;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= avisoRonda;
                    END IF;

                    letra3 <= '0';

                    letra2 <= '0';

                    letra1 <= '0';

                    letra0 <= '1';
                WHEN inputRonda =>
                    IF ((aceptar = '0')) THEN
                        reg_fstate <= ptosJugadores;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= inputRonda;
                    END IF;

                    letra3 <= '0';

                    letra2 <= '0';

                    letra1 <= '0';

                    letra0 <= '1';
						  
                WHEN ptosJugadores =>
                    IF ((aceptar = '1')) THEN
                        reg_fstate <= registroPtos;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ptosJugadores;
                    END IF;

                    letra3 <= '1';

                    letra2 <= '1';

                    letra1 <= '1';

                    letra0 <= '0';
                WHEN registroPtos =>
                    IF ((aceptar = '1')) THEN
                        reg_fstate <= inputPtos;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= registroPtos;
                    END IF;

                    Q0 <= '0';

                    Q1 <= '1';
                WHEN inputPtos =>
                    IF ((aceptar = '0')) THEN
                        reg_fstate <= ptosJugadores;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= inputPtos;
                    END IF;
                WHEN OTHERS => 
                    Q1 <= 'X';
                    Q0 <= 'X';
                    letra0 <= 'X';
                    letra1 <= 'X';
                    letra2 <= 'X';
                    letra3 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
